module simple_assign(
    input wire in,  // Input signal
    output wire out // Output signal
);
    // Assign the output to the input
    assign out = in;
endmodule
